module Mul_by2_Nbit #(parameter N = 8) (a,y);

input [N-1:0]a;
output [N-1:0]y;

assign y = {a[N-2:0],1'b0};

endmodule
