module Xnor_2in_Nbit #(parameter N = 8)(c,a,b);

input [N-1:0]a;
input [N-1:0]b;
output [N-1:0]c;

wire [N-1:0]a_bar;
wire [N-1:0]b_bar;
wire [N-1:0]y1;
wire [N-1:0]y2;
wire [N-1:0]y;

assign a_bar = ~a;
assign b_bar = ~b;
assign y1 = a&b_bar;
assign y2 = a_bar&b;
assign y = y1|y2;

assign c = ~y;

endmodule
