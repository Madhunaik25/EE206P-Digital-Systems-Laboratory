module TB_Top_assign1();

  parameter M = 4;

  reg [2:0]s;
  reg [M-1:0]a;
  reg [M-1:0]b;
  wire [M-1:0]c;

  Top_assign1 #(.N(M)) DUT(.a(a),.s(s),.b(b),.c(c));

  initial

  begin

/*    s = 3'b000; a = 4'b1001; b = 4'b1010;
    #10 
    s = 3'b001; a = 4'b0100; b = 4'b1000;
    #10
    s = 3'b010; a = 4'b1001; b = 4'b1010;
    #10
    s = 3'b011; a = 4'b0100; b = 4'b1000;
    #10
    s = 3'b100; a = 4'b1110; b = 4'b0111;
    #10
    s = 3'b101; a = 4'b1110; b = 4'b0111;
    #10
    s = 3'b110; a = 4'b0011; b = 4'b0000;
    #10
    s = 3'b111; a = 4'b0110; b = 4'b0000;
    #10;
*/
repeat(20)
begin
s = $random(); 
a = $random();
b = $random();
#10;
#5 $display("%b, %b, %b, %b", s, a, b, c );
end
$finish;   
end
initial



begin
$monitor("s = %b,a = %b,b = %b,c = %b", s, a, b, c );
end
endmodule 